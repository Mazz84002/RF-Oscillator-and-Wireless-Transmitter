** Profile: "SCHEMATIC1-bias-point"  [ c:\cadence_projects\final-design\collpits-oscillator-final-design-PSpiceFiles\SCHEMATIC1\bias-point.sim ] 

** Creating circuit file "bias-point.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\mazz\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.SAVEBIAS "C:/Cadence_Projects/Final-Design/Collpits-Oscillator-Final-Design-PSpiceFiles/SCHEMATIC1/bias-point/bias-point-output.txt" OP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
