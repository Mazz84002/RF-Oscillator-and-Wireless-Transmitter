** Profile: "SCHEMATIC1-ac-sweep"  [ C:\VCO-transmitter\Update-Oscillator-Design\Updated-Coll-pits-Oscillator-Design-PSpiceFiles\SCHEMATIC1\ac-sweep.sim ] 

** Creating circuit file "ac-sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\mazz\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC LIN 1000 1e9 5e9
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
