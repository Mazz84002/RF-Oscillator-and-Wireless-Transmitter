** Profile: "SCHEMATIC1-param-sweep"  [ C:\VCO-transmitter\PSpice-Load-Sweep\Load-sweep-PSpiceFiles\SCHEMATIC1\param-sweep.sim ] 

** Creating circuit file "param-sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\mazz\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 8e-8 0 1e-11 
.STEP LIN PARAM RL 540 1240 100 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
